/*
*Author : Revanth Sai Nandamuri
*GitHUB : https://github.com/RevanthNandamuri1341b0
*Date of update : 22 August 2021
*Project name : ALU Verification Environment
*Domain : UVM
*Description : Pre-defined Sequencer
*File Name : sequencer.sv
*File ID : 412157
*Modified by : #your name#
*/

typedef uvm_sequencer #(alu_trans) sequencer;